//===========================================================================
//-- File Version    : 1.00
//-- Date            : 25/11/25
//-- Author          : phong
//-- IP Name         : synchronizer 
//-- History         : ver.1.00 (25/11/24) 1st release
//--
//===========================================================================
module synchronizer #(
    parameter P_DATA_W = 8
)(
    input                               clk, 
    input                               rst_n, 
    input       [P_DATA_W - 1   : 0]    i_data, 
    output  reg [P_DATA_W - 1   : 0]    o_data
);
//---------------------------------------------------------------------------
    // PARAMETER HERE
//---------------------------------------------------------------------------
    // VARIABLE
    reg [P_DATA_W - 1   : 0]    q1;
//---------------------------------------------------------------------------
    always @(posedge clk) begin
        if(!rst_n) begin
            q1      <= 0;
            o_data  <= 0;
        end else begin
            q1      <= i_data;
            o_data  <= q1;
        end
    end
//---------------------------------------------------------------------------
endmodule
//===========================================================================