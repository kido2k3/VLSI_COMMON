//===========================================================================
//-- File Version    : 
//-- Date            : 
//-- Author          : kido
//-- All coverages are common in design verification, and its explaination
//===========================================================================
